module sum(
    input logic [19:0] n,  //Numero que esta entrando por el debounce
    output logic [9:0] s   //Suma de los 2 numeros
);


endmodule